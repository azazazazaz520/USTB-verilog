module top_module(
    input clk,
    input areset,    
    input in,
    output out
);
    
endmodule